"Test Save"

PLAYER_X
800

PLAYER_Y
800